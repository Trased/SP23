module ALU_tb;
reg [7:0] A;
reg [7:0] B;
reg [3:0] Sel;
wire [7:0] Out;
wire [3:0] Flag;

ALU alu_DUT(
            .A(A),
            .B(B),
            .Sel(Sel),
            .Out(Out),
            .Flag(Flag));
            
initial
begin
    #0
        A <= 8'h0;
        B <= 8'h0;
        Sel <= 4'h0;
    #10
        A <= 8'hC1;
        B <= 8'h0F;
    #10
        A <= 8'hFF;
        B <= 8'hFF;
    
    #10
        Sel <= 4'h1;
    #10
        A <= 8'hC1;
        B <= 8'h0F;
    #10
        A <= 8'h0F;
        B <= 8'hC1;       
    #10
        Sel <= 4'h2;
    #10
        A <= 8'hC1;
        B <= 8'h0F;
    #10
        A <= 8'h1F;
        B <= 8'h1F;
    #10
        Sel <= 4'h3;
    #10
        A <= 8'hC1;
        B <= 8'h0F;
    #10
        A <= 8'h0F;
        B <= 8'hC1;  
    #10
        Sel <= 4'h4;
        A <= 8'hFF;
        B <= 8'h4;
    #10
        B <= 8'h2;
    #10
        Sel <= 4'h5;
    #10
        B <= 8'h4;
    #10
        Sel <= 4'h6;
        A <= 8'b10101010;
        B <= 8'b10100000;
    #10
        B <= 8'b00000000;
    #10
        B <= 8'b11111111;
    #10
        Sel <= 4'h7;
    #10
        B <= 8'b01010101;
    #10
        A <= 8'b00001100;
        B <= 8'b11000011;
    #10
        Sel <= 4'h8;
        B <= 8'b10001111;
    #10
        A <= 8'b01110000;
    #10
        Sel <= 4'h9;
    #10
        B <= 8'b01010101;
    #10
        A <= 8'b00001100;
        B <= 8'b11000011;
    #10
        Sel <= 4'hA;
        A <= 8'b10101010;
        B <= 8'b10100000;
    #10
        B <= 8'b00000000;
    #10
        B <= 8'b11111111;
    #10
        Sel <= 4'hB;
    #10
        B <= 8'b01010101;
    #10
        A <= 8'b00001100;
        B <= 8'b11000011;
    #10
        Sel <= 4'hC;
    #10
        Sel <= 4'hE;    
    
        
    #10
        $finish;    
        
end

endmodule
